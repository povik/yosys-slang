module top;
initial begin
$t(1 + 1);
end
endmodule
