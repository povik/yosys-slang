module top;
	f f();
endmodule
