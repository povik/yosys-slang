`timescale 1ns/1ps

module f;
endmodule
